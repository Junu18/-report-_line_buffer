`include "line_buf_ctrl.v"
`include "top.v"
`include "single_port_ram.v"
