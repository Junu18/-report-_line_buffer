`include "top.v"
`include "single_port_ram.v"